module LZD #(parameter WIDTH = 25) (
    input logic [WIDTH-1:0] in, // in 
    output logic [$clog2(WIDTH):0] lead_zero_count // LZD count
);

    always_comb begin
        // Initialize the output to 0
        // Check from MSB to LSB, using a decoder-like structure
        casez (in)
            25'b1????????????????????????: lead_zero_count = 0;  // 
            25'b01???????????????????????: lead_zero_count = 1;  // 为1
            25'b001??????????????????????: lead_zero_count = 2;  // 
            25'b0001?????????????????????: lead_zero_count = 3;  // 
            25'b00001????????????????????: lead_zero_count = 4;  // 
            25'b000001???????????????????: lead_zero_count = 5;  // 
            25'b0000001??????????????????: lead_zero_count = 6;  // 
            25'b00000001?????????????????: lead_zero_count = 7;  // 
            25'b000000001????????????????: lead_zero_count = 8;  // 
            25'b0000000001???????????????: lead_zero_count = 9;  // 
            25'b00000000001??????????????: lead_zero_count = 10; // 
            25'b000000000001?????????????: lead_zero_count = 11; // 
            25'b0000000000001????????????: lead_zero_count = 12; // 
            25'b00000000000001???????????: lead_zero_count = 13; // 
            25'b000000000000001??????????: lead_zero_count = 14; // 
            25'b0000000000000001?????????: lead_zero_count = 15; // 
            25'b00000000000000001????????: lead_zero_count = 16; // 
            25'b000000000000000001???????: lead_zero_count = 17; // 
            25'b0000000000000000001??????: lead_zero_count = 18; // 
            25'b00000000000000000001?????: lead_zero_count = 19; // 
            25'b000000000000000000001????: lead_zero_count = 20; // 
            25'b0000000000000000000001???: lead_zero_count = 21; // 
            25'b00000000000000000000001??: lead_zero_count = 22; // 
            25'b000000000000000000000001?: lead_zero_count = 23; // 
            25'b0000000000000000000000001: lead_zero_count = 24; // 
            default: lead_zero_count = 25;                         // 
        endcase
    end

endmodule
