`define FLOAT_32_EXP 8
`define FLOAT_32_FRAC 23
`define ADD 1'b0
`define SUB 1'b1
`define FAR_PATH 1'b0
`define CLOSE_PATH 1'b1
`define Q_NaN 1'b1
`define S_NaN 1'b0