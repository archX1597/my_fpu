import FPU_pkg::*;
module FMA(
    input float_type OP_A,
    input float_type OP_B,
    input float_type OP_C
);

endmodule